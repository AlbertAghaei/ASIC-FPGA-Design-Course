module fft_radix2_16 (
    input wire clk,
    input wire rst,

    // Real and Imaginary inputs (16 complex numbers)
    input wire signed [15:0] real_in0,  input wire signed [15:0] imag_in0,
    input wire signed [15:0] real_in1,  input wire signed [15:0] imag_in1,
    input wire signed [15:0] real_in2,  input wire signed [15:0] imag_in2,
    input wire signed [15:0] real_in3,  input wire signed [15:0] imag_in3,
    input wire signed [15:0] real_in4,  input wire signed [15:0] imag_in4,
    input wire signed [15:0] real_in5,  input wire signed [15:0] imag_in5,
    input wire signed [15:0] real_in6,  input wire signed [15:0] imag_in6,
    input wire signed [15:0] real_in7,  input wire signed [15:0] imag_in7,
    input wire signed [15:0] real_in8,  input wire signed [15:0] imag_in8,
    input wire signed [15:0] real_in9,  input wire signed [15:0] imag_in9,
    input wire signed [15:0] real_in10, input wire signed [15:0] imag_in10,
    input wire signed [15:0] real_in11, input wire signed [15:0] imag_in11,
    input wire signed [15:0] real_in12, input wire signed [15:0] imag_in12,
    input wire signed [15:0] real_in13, input wire signed [15:0] imag_in13,
    input wire signed [15:0] real_in14, input wire signed [15:0] imag_in14,
    input wire signed [15:0] real_in15, input wire signed [15:0] imag_in15,

    // Real and Imaginary outputs
    output wire signed [15:0] real_out0,  output wire signed [15:0] imag_out0,
    output wire signed [15:0] real_out1,  output wire signed [15:0] imag_out1,
    output wire signed [15:0] real_out2,  output wire signed [15:0] imag_out2,
    output wire signed [15:0] real_out3,  output wire signed [15:0] imag_out3,
    output wire signed [15:0] real_out4,  output wire signed [15:0] imag_out4,
    output wire signed [15:0] real_out5,  output wire signed [15:0] imag_out5,
    output wire signed [15:0] real_out6,  output wire signed [15:0] imag_out6,
    output wire signed [15:0] real_out7,  output wire signed [15:0] imag_out7,
    output wire signed [15:0] real_out8,  output wire signed [15:0] imag_out8,
    output wire signed [15:0] real_out9,  output wire signed [15:0] imag_out9,
    output wire signed [15:0] real_out10, output wire signed [15:0] imag_out10,
    output wire signed [15:0] real_out11, output wire signed [15:0] imag_out11,
    output wire signed [15:0] real_out12, output wire signed [15:0] imag_out12,
    output wire signed [15:0] real_out13, output wire signed [15:0] imag_out13,
    output wire signed [15:0] real_out14, output wire signed [15:0] imag_out14,
    output wire signed [15:0] real_out15, output wire signed [15:0] imag_out15
);

   // Intermediate signals between stages
    wire signed [15:0] s1_r[15:0], s1_i[15:0];
    wire signed [15:0] s2_r[15:0], s2_i[15:0];
    wire signed [15:0] s3_r[15:0], s3_i[15:0];

    // Stage 1: First FFT layer
    fft_radix2_16_stage1 stage1 (
        .clk(clk), .rst(rst),
        .real_in0(real_in0), .imag_in0(imag_in0),
        .real_in1(real_in1), .imag_in1(imag_in1),
        .real_in2(real_in2), .imag_in2(imag_in2),
        .real_in3(real_in3), .imag_in3(imag_in3),
        .real_in4(real_in4), .imag_in4(imag_in4),
        .real_in5(real_in5), .imag_in5(imag_in5),
        .real_in6(real_in6), .imag_in6(imag_in6),
        .real_in7(real_in7), .imag_in7(imag_in7),
        .real_in8(real_in8), .imag_in8(imag_in8),
        .real_in9(real_in9), .imag_in9(imag_in9),
        .real_in10(real_in10), .imag_in10(imag_in10),
        .real_in11(real_in11), .imag_in11(imag_in11),
        .real_in12(real_in12), .imag_in12(imag_in12),
        .real_in13(real_in13), .imag_in13(imag_in13),
        .real_in14(real_in14), .imag_in14(imag_in14),
        .real_in15(real_in15), .imag_in15(imag_in15),
        .real_out0(s1_r[0]), .imag_out0(s1_i[0]),
        .real_out1(s1_r[1]), .imag_out1(s1_i[1]),
        .real_out2(s1_r[2]), .imag_out2(s1_i[2]),
        .real_out3(s1_r[3]), .imag_out3(s1_i[3]),
        .real_out4(s1_r[4]), .imag_out4(s1_i[4]),
        .real_out5(s1_r[5]), .imag_out5(s1_i[5]),
        .real_out6(s1_r[6]), .imag_out6(s1_i[6]),
        .real_out7(s1_r[7]), .imag_out7(s1_i[7]),
        .real_out8(s1_r[8]), .imag_out8(s1_i[8]),
        .real_out9(s1_r[9]), .imag_out9(s1_i[9]),
        .real_out10(s1_r[10]), .imag_out10(s1_i[10]),
        .real_out11(s1_r[11]), .imag_out11(s1_i[11]),
        .real_out12(s1_r[12]), .imag_out12(s1_i[12]),
        .real_out13(s1_r[13]), .imag_out13(s1_i[13]),
        .real_out14(s1_r[14]), .imag_out14(s1_i[14]),
        .real_out15(s1_r[15]), .imag_out15(s1_i[15])
    );

    // Stage 2: Twiddle W0, W2, W4, W6
    fft_radix2_16_stage2 stage2 (
        .clk(clk), .rst(rst),
        .real_in0(s1_r[0]), .imag_in0(s1_i[0]),
        .real_in1(s1_r[1]), .imag_in1(s1_i[1]),
        .real_in2(s1_r[2]), .imag_in2(s1_i[2]),
        .real_in3(s1_r[3]), .imag_in3(s1_i[3]),
        .real_in4(s1_r[4]), .imag_in4(s1_i[4]),
        .real_in5(s1_r[5]), .imag_in5(s1_i[5]),
        .real_in6(s1_r[6]), .imag_in6(s1_i[6]),
        .real_in7(s1_r[7]), .imag_in7(s1_i[7]),
        .real_in8(s1_r[8]), .imag_in8(s1_i[8]),
        .real_in9(s1_r[9]), .imag_in9(s1_i[9]),
        .real_in10(s1_r[10]), .imag_in10(s1_i[10]),
        .real_in11(s1_r[11]), .imag_in11(s1_i[11]),
        .real_in12(s1_r[12]), .imag_in12(s1_i[12]),
        .real_in13(s1_r[13]), .imag_in13(s1_i[13]),
        .real_in14(s1_r[14]), .imag_in14(s1_i[14]),
        .real_in15(s1_r[15]), .imag_in15(s1_i[15]),
        .real_out0(s2_r[0]), .imag_out0(s2_i[0]),
        .real_out1(s2_r[1]), .imag_out1(s2_i[1]),
        .real_out2(s2_r[2]), .imag_out2(s2_i[2]),
        .real_out3(s2_r[3]), .imag_out3(s2_i[3]),
        .real_out4(s2_r[4]), .imag_out4(s2_i[4]),
        .real_out5(s2_r[5]), .imag_out5(s2_i[5]),
        .real_out6(s2_r[6]), .imag_out6(s2_i[6]),
        .real_out7(s2_r[7]), .imag_out7(s2_i[7]),
        .real_out8(s2_r[8]), .imag_out8(s2_i[8]),
        .real_out9(s2_r[9]), .imag_out9(s2_i[9]),
        .real_out10(s2_r[10]), .imag_out10(s2_i[10]),
        .real_out11(s2_r[11]), .imag_out11(s2_i[11]),
        .real_out12(s2_r[12]), .imag_out12(s2_i[12]),
        .real_out13(s2_r[13]), .imag_out13(s2_i[13]),
        .real_out14(s2_r[14]), .imag_out14(s2_i[14]),
        .real_out15(s2_r[15]), .imag_out15(s2_i[15])
    );

    // Stage 3: Using only W = �1
    fft_radix2_16_stage3 stage3 (
        .clk(clk), .rst(rst),
        .real_in0(s2_r[0]), .imag_in0(s2_i[0]),
        .real_in1(s2_r[1]), .imag_in1(s2_i[1]),
        .real_in2(s2_r[2]), .imag_in2(s2_i[2]),
        .real_in3(s2_r[3]), .imag_in3(s2_i[3]),
        .real_in4(s2_r[4]), .imag_in4(s2_i[4]),
        .real_in5(s2_r[5]), .imag_in5(s2_i[5]),
        .real_in6(s2_r[6]), .imag_in6(s2_i[6]),
        .real_in7(s2_r[7]), .imag_in7(s2_i[7]),
        .real_in8(s2_r[8]), .imag_in8(s2_i[8]),
        .real_in9(s2_r[9]), .imag_in9(s2_i[9]),
        .real_in10(s2_r[10]), .imag_in10(s2_i[10]),
        .real_in11(s2_r[11]), .imag_in11(s2_i[11]),
        .real_in12(s2_r[12]), .imag_in12(s2_i[12]),
        .real_in13(s2_r[13]), .imag_in13(s2_i[13]),
        .real_in14(s2_r[14]), .imag_in14(s2_i[14]),
        .real_in15(s2_r[15]), .imag_in15(s2_i[15]),
        .real_out0(s3_r[0]), .imag_out0(s3_i[0]),
        .real_out1(s3_r[1]), .imag_out1(s3_i[1]),
        .real_out2(s3_r[2]), .imag_out2(s3_i[2]),
        .real_out3(s3_r[3]), .imag_out3(s3_i[3]),
        .real_out4(s3_r[4]), .imag_out4(s3_i[4]),
        .real_out5(s3_r[5]), .imag_out5(s3_i[5]),
        .real_out6(s3_r[6]), .imag_out6(s3_i[6]),
        .real_out7(s3_r[7]), .imag_out7(s3_i[7]),
        .real_out8(s3_r[8]), .imag_out8(s3_i[8]),
        .real_out9(s3_r[9]), .imag_out9(s3_i[9]),
        .real_out10(s3_r[10]), .imag_out10(s3_i[10]),
        .real_out11(s3_r[11]), .imag_out11(s3_i[11]),
        .real_out12(s3_r[12]), .imag_out12(s3_i[12]),
        .real_out13(s3_r[13]), .imag_out13(s3_i[13]),
        .real_out14(s3_r[14]), .imag_out14(s3_i[14]),
        .real_out15(s3_r[15]), .imag_out15(s3_i[15])
    );

    // Stage 4: Final summation stage (no twiddle)
    fft_radix2_16_stage4 stage4 (
        .clk(clk), .rst(rst),
        .real_in0(s3_r[0]), .imag_in0(s3_i[0]),
        .real_in1(s3_r[1]), .imag_in1(s3_i[1]),
        .real_in2(s3_r[2]), .imag_in2(s3_i[2]),
        .real_in3(s3_r[3]), .imag_in3(s3_i[3]),
        .real_in4(s3_r[4]), .imag_in4(s3_i[4]),
        .real_in5(s3_r[5]), .imag_in5(s3_i[5]),
        .real_in6(s3_r[6]), .imag_in6(s3_i[6]),
        .real_in7(s3_r[7]), .imag_in7(s3_i[7]),
        .real_in8(s3_r[8]), .imag_in8(s3_i[8]),
        .real_in9(s3_r[9]), .imag_in9(s3_i[9]),
        .real_in10(s3_r[10]), .imag_in10(s3_i[10]),
        .real_in11(s3_r[11]), .imag_in11(s3_i[11]),
        .real_in12(s3_r[12]), .imag_in12(s3_i[12]),
        .real_in13(s3_r[13]), .imag_in13(s3_i[13]),
        .real_in14(s3_r[14]), .imag_in14(s3_i[14]),
        .real_in15(s3_r[15]), .imag_in15(s3_i[15]),
        .real_out0(real_out0),   .imag_out0(imag_out0),
        .real_out1(real_out1),   .imag_out1(imag_out1),
        .real_out2(real_out2),   .imag_out2(imag_out2),
        .real_out3(real_out3),   .imag_out3(imag_out3),
        .real_out4(real_out4),   .imag_out4(imag_out4),
        .real_out5(real_out5),   .imag_out5(imag_out5),
        .real_out6(real_out6),   .imag_out6(imag_out6),
        .real_out7(real_out7),   .imag_out7(imag_out7),
        .real_out8(real_out8),   .imag_out8(imag_out8),
        .real_out9(real_out9),   .imag_out9(imag_out9),
        .real_out10(real_out10), .imag_out10(imag_out10),
        .real_out11(real_out11), .imag_out11(imag_out11),
        .real_out12(real_out12), .imag_out12(imag_out12),
        .real_out13(real_out13), .imag_out13(imag_out13),
        .real_out14(real_out14), .imag_out14(imag_out14),
        .real_out15(real_out15), .imag_out15(imag_out15)
    );

endmodule
